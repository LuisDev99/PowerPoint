// VGA protocol constants for 800x600 resolution
`define VGA_WIDTH  800
`define VGA_HEIGHT 600
`define VGA_HLIMIT 1056
`define VGA_VLIMIT 628
`define VGA_HSYNC_PULSE_START 840
`define VGA_HSYNC_PULSE_END   968
`define VGA_VSYNC_PULSE_START 601
`define VGA_VSYNC_PULSE_END   605

`define COLOR_BITS 8